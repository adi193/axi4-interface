package axi_stream_pkg;

	localparam DATA_WIDTH = 32;

	typedef logic [DATA_WIDTH - 1 : 0] data_t;

endpackage
